
module top(
	input wire clk
);
	initial begin
		$display("This is, a MESSAGE.");
	end
endmodule
